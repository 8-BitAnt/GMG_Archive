  S L           ����      Y@�   �	     �    ��            @        ��           �?        ��                     ��                     ��            @        ��           �?        ��                     ��           �?        ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                                          Æ                     Ć                     ņ                     Ɔ                     ǆ                     Ȇ                     Ɇ                     ʆ                     ˆ                     ̆                     ͆                     Ά                     φ                     І                     ц                     ҆                     ӆ                     Ԇ                     Ն                     ֆ                     ׆           �?        ؆                     ن          �@        چ                     ۆ                     ܆           b@        ݆           e@        ކ                     ߆                     ��           �?        �                     �                     �                     �                     �           �?        �                     �            @        �           @        �            @        Ȉ           �?        Ɉ                     ��               file    ƈ           @        ň           �?        ʈ           �?        ��                     ��                     ˈ            @        �         @[�@        Έ         @v�@        ͈           �?        ��                     ��            	   Your name    ��               Name of your level    ��           �?        ̈                     ψ               customlevelx.lef    �            @        �            @        �            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @         �            @        �            @        �            @        �            @        �            @        �            @        �            @        �            @        �            @        	�            @        
�            @        �            @        �            @        �            @        �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                      �                     !�                     "�                     #�                     $�                     %�                     &�                     '�            @        (�            @        )�                     *�                     +�                     ,�                     -�                     .�                     /�                     0�                     1�                     2�                     3�                     4�                     5�                     6�                     7�                     8�                     9�                     :�                     ;�                     <�                     =�                     >�                     ?�                     @�                     A�                     B�            @        C�            @        D�                     E�                     F�                     G�                     H�                     I�                     J�                     K�                     L�                     M�                     N�                     O�                     P�                     Q�                     R�                     S�                     T�                     U�                     V�                     W�                     X�                     Y�                     Z�                     [�                     \�                     ]�            @        ^�            @        _�                     `�                     a�                     b�                     c�                     d�                     e�                     f�                     g�                     h�                     i�                     j�                     k�                     l�                     m�                     n�                     o�                     p�                     q�                     r�                     s�                     t�                     u�                     v�                     w�                     x�            @        y�            @        z�                     {�                     |�                     }�                     ~�                     �                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��            @        ��            @        ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��            @        ��            @        ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                                          Ç                     ć                     Ň                     Ƈ                     Ǉ                     ȇ                     ɇ            @        ʇ            @        ˇ                     ̇                     ͇                     ·                     χ                     Ї                     ч                     ҇                     Ӈ                     ԇ                     Շ                     և                     ׇ                     ؇                     ه                     ڇ                     ۇ                     ܇                     ݇                     އ                     ߇                     ��                     �                     �                     �                     �            @        �            @        �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     ��                     �                     �                     �                     �                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��                     ��            @         �            @        �                     �                     �                     �                     �                     �                     �                     �                     	�                     
�                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �            @        �            @        �                     �                     �                     �                      �                     !�                     "�                     #�                     $�                     %�                     &�                     '�                     (�                     )�                     *�                     +�                     ,�                     -�                     .�                     /�                     0�                     1�                     2�                     3�                     4�                     5�            @        6�            @        7�                     8�                     9�                     :�                     ;�                     <�                     =�                     >�                     ?�                     @�                     A�                     B�                     C�                     D�                     E�                     F�                     G�                     H�                     I�                     J�                     K�                     L�                     M�                     N�                     O�                     P�            @        Q�            @        R�                     S�                     T�                     U�                     V�                     W�                     X�                     Y�                     Z�                     [�                     \�                     ]�                     ^�                     _�                     `�                     a�                     b�                     c�                     d�                     e�                     f�                     g�                     h�                     i�                     j�                     k�            @        l�            @        m�                     n�                     o�                     p�                     q�                     r�                     s�                     t�                     u�                     v�                     w�                     x�                     y�                     z�                     {�                     |�                     }�                     ~�                     �                     ��                     ��                     ��                     ��                     ��                     ��                     ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        ��            @        "                                                                                                                                                                                                                                                                                                                           �  �  <              q   script_levelstart()

instance_create(0,0,mouse_on)

if file_exists("basic.lef")
{
game_load("basic.lef")
}                                          �?      �?                ���       �?        ����                            �?      �?                ���       �?        ����                            �?      �?                ���       �?        ����                            �?      �?                ���       �?        ����                            �?      �?                ���       �?        ����                            �?      �?                ���       �?        ����                            �?      �?                ���       �?        ����                            �?      �?                ���       �?                   �  �          �  �                  ������������            �  �          �  �                  ������������            �  �          �  �                  ������������            �  �          �  �                  ������������            �  �          �  �                  ������������            �  �          �  �                  ������������            �  �          �  �                  ������������            �  �          �  �                  ������������  �� ����     X�@      �?      �?      �?              �?��� ����                                                                                         �p@                        `y��`y��`y��`y��           �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t          @              �?      �?              �?��� ����                         {@              {@              {@                             �p@                               �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t          @              �?      �?              �?���                              H@              H@              H@                             �p@                               0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           �?        ��                     �� t          @              �?      �?              �?���                      8@      H@      8@      H@      8@      H@                             �p@                           /   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��            @        ��                     �� t          @              �?      �?              �?���                      H@      H@      H@      H@      H@      H@                             �p@                        0   G   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           @        ��                     �� t          @              �?      �?              �?���                      R@      H@      R@      H@      R@      H@                             �p@                        H   _   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           @        ��                     �� t          @              �?      �?              �?���                      X@      H@      X@      H@      X@      H@                             �p@                        `   w   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           @        ��                     �� t          @              �?      �?              �?���                      ^@      H@      ^@      H@      ^@      H@                             �p@                        x   �   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           @        ��                     �� t          @              �?      �?              �?���                      b@      H@      b@      H@      b@      H@                             �p@                        �   �   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           @        ��                     �� t          @              �?      �?              �?���                      e@      H@      e@      H@      e@      H@                             �p@                        �   �   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��            @        ��                     �� t          @              �?      �?              �?���                      h@      H@      h@      H@      h@      H@                             �p@                        �   �   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           "@        ��                     �� t          @              �?      �?              �?���                      k@      H@      k@      H@      k@      H@                             �p@                        �   �   0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           $@        ��                     �� t          @              �?      �?              �?���                      n@      H@      n@      H@      n@      H@                             �p@                        �     0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           &@        ��                     �� t          @              �?      �?              �?���                     �p@      H@     �p@      H@     �p@      H@                             �p@                            0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           (@        ��                     �� t          @              �?      �?              �?���                      r@      H@      r@      H@      r@      H@                             �p@                           7  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           *@        ��                     �� t          @              �?      �?              �?���                     �s@      H@     �s@      H@     �s@      H@                             �p@                        8  O  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           ,@        ��                     �� t          @              �?      �?              �?���                      u@      H@      u@      H@      u@      H@                             �p@                        P  g  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           .@        ��                     �� t          @              �?      �?              �?���                     �v@      H@     �v@      H@     �v@      H@                             �p@                        h    0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           0@        ��                     �� t          @              �?      �?              �?���                      x@      H@      x@      H@      x@      H@                             �p@                        �  �  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           1@        ��                     �� t          @              �?      �?              �?���                     �y@      H@     �y@      H@     �y@      H@                             �p@                        �  �  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           2@        ��                     �� t          @              �?      �?              �?���                      {@      H@      {@      H@      {@      H@                             �p@                        �  �  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           3@        ��                     �� t          @              �?      �?              �?���                     �|@      H@     �|@      H@     �|@      H@                             �p@                        �  �  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           4@        ��                     �� t          @              �?      �?              �?���                      ~@      H@      ~@      H@      ~@      H@                             �p@                        �  �  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           5@        ��                     �� t          @              �?      �?              �?���                     �@      H@     �@      H@     �@      H@                             �p@                        �    0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           6@        ��                     �� t          @              �?      �?              �?���                     ��@      H@     ��@      H@     ��@      H@                             �p@                          '  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           7@        ��                     �� t          @              �?      �?              �?���                     @�@      H@     @�@      H@     @�@      H@                             �p@                        (  ?  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           8@        ��                     �� t          @              �?      �?              �?���                      �@      H@      �@      H@      �@      H@                             �p@                        @  W  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           9@        ��                     �� t          @              �?      �?              �?���                     ��@      H@     ��@      H@     ��@      H@                             �p@                        X  o  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           :@        ��                     �� t          @              �?      �?              �?���                     ��@      H@     ��@      H@     ��@      H@                             �p@                        p  �  0   G              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           ;@        ��                     �� t          @              �?      �?              �?���                              R@              R@              R@                             �p@                               H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           <@        ��                     �� t                         �?      �?              �?���                      8@      R@      8@      R@      8@      R@                             �p@                           /   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           =@        ��                     �� t                         �?      �?              �?���                      H@      R@      H@      R@      H@      R@                             �p@                        0   G   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           >@        ��                     �� t                         �?      �?              �?���                      R@      R@      R@      R@      R@      R@                             �p@                        H   _   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           ?@        ��                     �� t                         �?      �?              �?���                      X@      R@      X@      R@      X@      R@                             �p@                        `   w   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           @@        ��                     �� t                         �?      �?              �?���                      ^@      R@      ^@      R@      ^@      R@                             �p@                        x   �   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �@@        ��                     �� t                         �?      �?              �?���                      b@      R@      b@      R@      b@      R@                             �p@                        �   �   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           A@        ��                     �� t                         �?      �?              �?���                      e@      R@      e@      R@      e@      R@                             �p@                        �   �   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �A@        ��                     �� t                         �?      �?              �?���                      h@      R@      h@      R@      h@      R@                             �p@                        �   �   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           B@        ��                     �� t                         �?      �?              �?���                      k@      R@      k@      R@      k@      R@                             �p@                        �   �   H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �B@        ��                     �� t                         �?      �?              �?���                      n@      R@      n@      R@      n@      R@                             �p@                        �     H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           C@        ��                     �� t                         �?      �?              �?���                     �p@      R@     �p@      R@     �p@      R@                             �p@                            H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �C@        ��                     �� t                         �?      �?              �?���                      r@      R@      r@      R@      r@      R@                             �p@                           7  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           D@        ��                     �� t                         �?      �?              �?���                     �s@      R@     �s@      R@     �s@      R@                             �p@                        8  O  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �D@        ��                     �� t                         �?      �?              �?���                      u@      R@      u@      R@      u@      R@                             �p@                        P  g  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           E@        ��                     �� t                         �?      �?              �?���                     �v@      R@     �v@      R@     �v@      R@                             �p@                        h    H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �E@        ��                     �� t                         �?      �?              �?���                      x@      R@      x@      R@      x@      R@                             �p@                        �  �  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           F@        ��                     �� t                         �?      �?              �?���                     �y@      R@     �y@      R@     �y@      R@                             �p@                        �  �  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �F@        ��                     �� t                         �?      �?              �?���                      {@      R@      {@      R@      {@      R@                             �p@                        �  �  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           G@        ��                     �� t                         �?      �?              �?���                     �|@      R@     �|@      R@     �|@      R@                             �p@                        �  �  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �G@        ��                     �� t                         �?      �?              �?���                      ~@      R@      ~@      R@      ~@      R@                             �p@                        �  �  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           H@        ��                     �� t                         �?      �?              �?���                     �@      R@     �@      R@     �@      R@                             �p@                        �    H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �H@        ��                     �� t                         �?      �?              �?���                     ��@      R@     ��@      R@     ��@      R@                             �p@                          '  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           I@        ��                     �� t                         �?      �?              �?���                     @�@      R@     @�@      R@     @�@      R@                             �p@                        (  ?  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �I@        ��                     �� t                         �?      �?              �?���                      �@      R@      �@      R@      �@      R@                             �p@                        @  W  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           J@        ��                     �� t                         �?      �?              �?���                     ��@      R@     ��@      R@     ��@      R@                             �p@                        X  o  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �J@        ��                     �� t          @              �?      �?              �?���                     ��@      R@     ��@      R@     ��@      R@                             �p@                        p  �  H   _              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           K@        ��                     �� t          @              �?      �?              �?���                              X@              X@              X@                             �p@                               `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �K@        ��                     �� t                         �?      �?              �?���                      8@      X@      8@      X@      8@      X@                             �p@                           /   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           L@        ��                     �� t                         �?      �?              �?���                      H@      X@      H@      X@      H@      X@                             �p@                        0   G   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �L@        ��                     �� t                         �?      �?              �?���                      R@      X@      R@      X@      R@      X@                             �p@                        H   _   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           M@        ��                     �� t                         �?      �?              �?���                      X@      X@      X@      X@      X@      X@                             �p@                        `   w   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �M@        ��                     �� t                         �?      �?              �?���                      ^@      X@      ^@      X@      ^@      X@                             �p@                        x   �   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           N@        ��                     �� t                         �?      �?              �?���                      b@      X@      b@      X@      b@      X@                             �p@                        �   �   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �N@        ��                     �� t                         �?      �?              �?���                      e@      X@      e@      X@      e@      X@                             �p@                        �   �   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           O@        ��                     �� t                         �?      �?              �?���                      h@      X@      h@      X@      h@      X@                             �p@                        �   �   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �O@        ��                     �� t                         �?      �?              �?���                      k@      X@      k@      X@      k@      X@                             �p@                        �   �   `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           P@        ��                     �� t                         �?      �?              �?���                      n@      X@      n@      X@      n@      X@                             �p@                        �     `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @P@        ��                     �� t                         �?      �?              �?���                     �p@      X@     �p@      X@     �p@      X@                             �p@                            `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �P@        ��                     �� t                         �?      �?              �?���                      r@      X@      r@      X@      r@      X@                             �p@                           7  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �P@        ��                     �� t                         �?      �?              �?���                     �s@      X@     �s@      X@     �s@      X@                             �p@                        8  O  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           Q@        ��                     �� t                         �?      �?              �?���                      u@      X@      u@      X@      u@      X@                             �p@                        P  g  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @Q@        ��                     �� t                         �?      �?              �?���                     �v@      X@     �v@      X@     �v@      X@                             �p@                        h    `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �Q@        ��                     �� t                         �?      �?              �?���                      x@      X@      x@      X@      x@      X@                             �p@                        �  �  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �Q@        ��                     �� t                         �?      �?              �?���                     �y@      X@     �y@      X@     �y@      X@                             �p@                        �  �  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           R@        ��                     �� t                         �?      �?              �?���                      {@      X@      {@      X@      {@      X@                             �p@                        �  �  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @R@        ��                     �� t                         �?      �?              �?���                     �|@      X@     �|@      X@     �|@      X@                             �p@                        �  �  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �R@        ��                     �� t                         �?      �?              �?���                      ~@      X@      ~@      X@      ~@      X@                             �p@                        �  �  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �R@        ��                     �� t                         �?      �?              �?���                     �@      X@     �@      X@     �@      X@                             �p@                        �    `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           S@        ��                      � t                         �?      �?              �?���                     ��@      X@     ��@      X@     ��@      X@                             �p@                          '  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @S@        ��                     � t                         �?      �?              �?���                     @�@      X@     @�@      X@     @�@      X@                             �p@                        (  ?  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �S@        ��                     � t                         �?      �?              �?���                      �@      X@      �@      X@      �@      X@                             �p@                        @  W  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �S@        ��                     � t                         �?      �?              �?���                     ��@      X@     ��@      X@     ��@      X@                             �p@                        X  o  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           T@        ��                     � t          @              �?      �?              �?���                     ��@      X@     ��@      X@     ��@      X@                             �p@                        p  �  `   w              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @T@        ��                     � t          @              �?      �?              �?���                              ^@              ^@              ^@                             �p@                               x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �T@        ��                     � t                         �?      �?              �?���                      8@      ^@      8@      ^@      8@      ^@                             �p@                           /   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �T@        ��                     � t                         �?      �?              �?���                      H@      ^@      H@      ^@      H@      ^@                             �p@                        0   G   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           U@        ��                     � t                         �?      �?              �?���                      R@      ^@      R@      ^@      R@      ^@                             �p@                        H   _   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @U@        ��                     	� t                         �?      �?              �?���                      X@      ^@      X@      ^@      X@      ^@                             �p@                        `   w   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �U@        ��                     
� t                         �?      �?              �?���                      ^@      ^@      ^@      ^@      ^@      ^@                             �p@                        x   �   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �U@        ��                     � t                         �?      �?              �?���                      b@      ^@      b@      ^@      b@      ^@                             �p@                        �   �   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           V@        ��                     � t                         �?      �?              �?���                      e@      ^@      e@      ^@      e@      ^@                             �p@                        �   �   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @V@        ��                     � t                         �?      �?              �?���                      h@      ^@      h@      ^@      h@      ^@                             �p@                        �   �   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �V@        ��                     � t                         �?      �?              �?���                      k@      ^@      k@      ^@      k@      ^@                             �p@                        �   �   x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �V@        ��                     � t                         �?      �?              �?���                      n@      ^@      n@      ^@      n@      ^@                             �p@                        �     x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           W@        ��                     � t                         �?      �?              �?���                     �p@      ^@     �p@      ^@     �p@      ^@                             �p@                            x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @W@        ��                     � t                         �?      �?              �?���                      r@      ^@      r@      ^@      r@      ^@                             �p@                           7  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �W@        ��                     � t                         �?      �?              �?���                     �s@      ^@     �s@      ^@     �s@      ^@                             �p@                        8  O  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �W@        ��                     � t                         �?      �?              �?���                      u@      ^@      u@      ^@      u@      ^@                             �p@                        P  g  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           X@        ��                     � t                         �?      �?              �?���                     �v@      ^@     �v@      ^@     �v@      ^@                             �p@                        h    x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @X@        ��                     � t                         �?      �?              �?���                      x@      ^@      x@      ^@      x@      ^@                             �p@                        �  �  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �X@        ��                     � t                         �?      �?              �?���                     �y@      ^@     �y@      ^@     �y@      ^@                             �p@                        �  �  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �X@        ��                     � t                         �?      �?              �?���                      {@      ^@      {@      ^@      {@      ^@                             �p@                        �  �  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           Y@        ��                     � t                         �?      �?              �?���                     �|@      ^@     �|@      ^@     �|@      ^@                             �p@                        �  �  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @Y@        ��                     � t                         �?      �?              �?���                      ~@      ^@      ~@      ^@      ~@      ^@                             �p@                        �  �  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �Y@        ��                     � t                         �?      �?              �?���                     �@      ^@     �@      ^@     �@      ^@                             �p@                        �    x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �Y@        ��                     � t                         �?      �?              �?���                     ��@      ^@     ��@      ^@     ��@      ^@                             �p@                          '  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           Z@        ��                     � t                         �?      �?              �?���                     @�@      ^@     @�@      ^@     @�@      ^@                             �p@                        (  ?  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @Z@        ��                     � t                         �?      �?              �?���                      �@      ^@      �@      ^@      �@      ^@                             �p@                        @  W  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �Z@        ��                     � t                         �?      �?              �?���                     ��@      ^@     ��@      ^@     ��@      ^@                             �p@                        X  o  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �Z@        ��                     � t          @              �?      �?              �?���                     ��@      ^@     ��@      ^@     ��@      ^@                             �p@                        p  �  x   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           [@        ��                      � t          @              �?      �?              �?���                              b@              b@              b@                             �p@                               �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @[@        ��                     !� t                         �?      �?              �?���                      8@      b@      8@      b@      8@      b@                             �p@                           /   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �[@        ��                     "� t                         �?      �?              �?���                      H@      b@      H@      b@      H@      b@                             �p@                        0   G   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �[@        ��                     #� t                         �?      �?              �?���                      R@      b@      R@      b@      R@      b@                             �p@                        H   _   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           \@        ��                     $� t                         �?      �?              �?���                      X@      b@      X@      b@      X@      b@                             �p@                        `   w   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @\@        ��                     %� t                         �?      �?              �?���                      ^@      b@      ^@      b@      ^@      b@                             �p@                        x   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �\@        ��                     &� t                         �?      �?              �?���                      b@      b@      b@      b@      b@      b@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �\@        ��                     '� t                         �?      �?              �?���                      e@      b@      e@      b@      e@      b@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           ]@        ��                     (� t                         �?      �?              �?���                      h@      b@      h@      b@      h@      b@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @]@        ��                     )� t                         �?      �?              �?���                      k@      b@      k@      b@      k@      b@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �]@        ��                     *� t                         �?      �?              �?���                      n@      b@      n@      b@      n@      b@                             �p@                        �     �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �]@        ��                     +� t                         �?      �?              �?���                     �p@      b@     �p@      b@     �p@      b@                             �p@                            �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           ^@        ��                     ,� t                         �?      �?              �?���                      r@      b@      r@      b@      r@      b@                             �p@                           7  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @^@        ��                     -� t                         �?      �?              �?���                     �s@      b@     �s@      b@     �s@      b@                             �p@                        8  O  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �^@        ��                     .� t                         �?      �?              �?���                      u@      b@      u@      b@      u@      b@                             �p@                        P  g  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �^@        ��                     /� t                         �?      �?              �?���                     �v@      b@     �v@      b@     �v@      b@                             �p@                        h    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           _@        ��                     0� t                         �?      �?              �?���                      x@      b@      x@      b@      x@      b@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @_@        ��                     1� t                         �?      �?              �?���                     �y@      b@     �y@      b@     �y@      b@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �_@        ��                     2� t                         �?      �?              �?���                      {@      b@      {@      b@      {@      b@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �_@        ��                     3� t                         �?      �?              �?���                     �|@      b@     �|@      b@     �|@      b@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           `@        ��                     4� t                         �?      �?              �?���                      ~@      b@      ~@      b@      ~@      b@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           `@        ��                     5� t                         �?      �?              �?���                     �@      b@     �@      b@     �@      b@                             �p@                        �    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @`@        ��                     6� t                         �?      �?              �?���                     ��@      b@     ��@      b@     ��@      b@                             �p@                          '  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          ``@        ��                     7� t                         �?      �?              �?���                     @�@      b@     @�@      b@     @�@      b@                             �p@                        (  ?  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �`@        ��                     8� t                         �?      �?              �?���                      �@      b@      �@      b@      �@      b@                             �p@                        @  W  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �`@        ��                     9� t                         �?      �?              �?���                     ��@      b@     ��@      b@     ��@      b@                             �p@                        X  o  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �`@        ��                     :� t          @              �?      �?              �?���                     ��@      b@     ��@      b@     ��@      b@                             �p@                        p  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �`@        ��                     ;� t          @              �?      �?              �?���                              e@              e@              e@                             �p@                               �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           a@        ��                     <� t                         �?      �?              �?���                      8@      e@      8@      e@      8@      e@                             �p@                           /   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           a@        ��                     =� t                         �?      �?              �?���                      H@      e@      H@      e@      H@      e@                             �p@                        0   G   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @a@        ��                     >� t                         �?      �?              �?���                      R@      e@      R@      e@      R@      e@                             �p@                        H   _   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `a@        ��                     ?� t                         �?      �?              �?���                      X@      e@      X@      e@      X@      e@                             �p@                        `   w   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �a@        ��                     @� t                         �?      �?              �?���                      ^@      e@      ^@      e@      ^@      e@                             �p@                        x   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �a@        ��                     A� t                         �?      �?              �?���                      b@      e@      b@      e@      b@      e@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �a@        ��                     B� t                         �?      �?              �?���                      e@      e@      e@      e@      e@      e@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �a@        ��                     C� t                         �?      �?              �?���                      h@      e@      h@      e@      h@      e@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           b@        ��                     D� t                         �?      �?              �?���                      k@      e@      k@      e@      k@      e@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           b@        ��                     E� t                         �?      �?              �?���                      n@      e@      n@      e@      n@      e@                             �p@                        �     �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @b@        ��                     F� t                         �?      �?              �?���                     �p@      e@     �p@      e@     �p@      e@                             �p@                            �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `b@        ��                     G� t                         �?      �?              �?���                      r@      e@      r@      e@      r@      e@                             �p@                           7  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �b@        ��                     H� t                         �?      �?              �?���                     �s@      e@     �s@      e@     �s@      e@                             �p@                        8  O  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �b@        ��                     I� t                         �?      �?              �?���                      u@      e@      u@      e@      u@      e@                             �p@                        P  g  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �b@        ��                     J� t                         �?      �?              �?���                     �v@      e@     �v@      e@     �v@      e@                             �p@                        h    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �b@        ��                     K� t                         �?      �?              �?���                      x@      e@      x@      e@      x@      e@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           c@        ��                     L� t                         �?      �?              �?���                     �y@      e@     �y@      e@     �y@      e@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           c@        ��                     M� t                         �?      �?              �?���                      {@      e@      {@      e@      {@      e@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @c@        ��                     N� t                         �?      �?              �?���                     �|@      e@     �|@      e@     �|@      e@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `c@        ��                     O� t                         �?      �?              �?���                      ~@      e@      ~@      e@      ~@      e@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �c@        ��                     P� t                         �?      �?              �?���                     �@      e@     �@      e@     �@      e@                             �p@                        �    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �c@        ��                     Q� t                         �?      �?              �?���                     ��@      e@     ��@      e@     ��@      e@                             �p@                          '  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �c@        ��                     R� t                         �?      �?              �?���                     @�@      e@     @�@      e@     @�@      e@                             �p@                        (  ?  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �c@        ��                     S� t                         �?      �?              �?���                      �@      e@      �@      e@      �@      e@                             �p@                        @  W  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           d@        ��                     T� t                         �?      �?              �?���                     ��@      e@     ��@      e@     ��@      e@                             �p@                        X  o  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           d@        ��                     U� t          @              �?      �?              �?���                     ��@      e@     ��@      e@     ��@      e@                             �p@                        p  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @d@        ��                     V� t          @              �?      �?              �?���                              h@              h@              h@                             �p@                               �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `d@        ��                     W� t                         �?      �?              �?���                      8@      h@      8@      h@      8@      h@                             �p@                           /   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �d@        ��                     X� t                         �?      �?              �?���                      H@      h@      H@      h@      H@      h@                             �p@                        0   G   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �d@        ��                     Y� t                         �?      �?              �?���                      R@      h@      R@      h@      R@      h@                             �p@                        H   _   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �d@        ��                     Z� t                         �?      �?              �?���                      X@      h@      X@      h@      X@      h@                             �p@                        `   w   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �d@        ��                     [� t                         �?      �?              �?���                      ^@      h@      ^@      h@      ^@      h@                             �p@                        x   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           e@        ��                     \� t                         �?      �?              �?���                      b@      h@      b@      h@      b@      h@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           e@        ��                     ]� t                         �?      �?              �?���                      e@      h@      e@      h@      e@      h@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @e@        ��                     ^� t                         �?      �?              �?���                      h@      h@      h@      h@      h@      h@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `e@        ��                     _� t                         �?      �?              �?���                      k@      h@      k@      h@      k@      h@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �e@        ��                     `� t                         �?      �?              �?���                      n@      h@      n@      h@      n@      h@                             �p@                        �     �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �e@        ��                     a� t                         �?      �?              �?���                     �p@      h@     �p@      h@     �p@      h@                             �p@                            �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �e@        ��                     b� t                         �?      �?              �?���                      r@      h@      r@      h@      r@      h@                             �p@                           7  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �e@        ��                     c� t                         �?      �?              �?���                     �s@      h@     �s@      h@     �s@      h@                             �p@                        8  O  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           f@        ��                     d� t                         �?      �?              �?���                      u@      h@      u@      h@      u@      h@                             �p@                        P  g  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           f@        ��                     e� t                         �?      �?              �?���                     �v@      h@     �v@      h@     �v@      h@                             �p@                        h    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @f@        ��                     f� t                         �?      �?              �?���                      x@      h@      x@      h@      x@      h@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `f@        ��                     g� t                         �?      �?              �?���                     �y@      h@     �y@      h@     �y@      h@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �f@        ��                     h� t                         �?      �?              �?���                      {@      h@      {@      h@      {@      h@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �f@        ��                     i� t                         �?      �?              �?���                     �|@      h@     �|@      h@     �|@      h@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �f@        ��                     j� t                         �?      �?              �?���                      ~@      h@      ~@      h@      ~@      h@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �f@        ��                     k� t                         �?      �?              �?���                     �@      h@     �@      h@     �@      h@                             �p@                        �    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           g@        ��                     l� t                         �?      �?              �?���                     ��@      h@     ��@      h@     ��@      h@                             �p@                          '  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           g@        ��                     m� t                         �?      �?              �?���                     @�@      h@     @�@      h@     @�@      h@                             �p@                        (  ?  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @g@        ��                     n� t                         �?      �?              �?���                      �@      h@      �@      h@      �@      h@                             �p@                        @  W  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `g@        ��                     o� t                         �?      �?              �?���                     ��@      h@     ��@      h@     ��@      h@                             �p@                        X  o  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �g@        ��                     p� t          @              �?      �?              �?���                     ��@      h@     ��@      h@     ��@      h@                             �p@                        p  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �g@        ��                     q� t          @              �?      �?              �?���                              k@              k@              k@                             �p@                               �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �g@        ��                     r� t                         �?      �?              �?���                      8@      k@      8@      k@      8@      k@                             �p@                           /   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �g@        ��                     s� t                         �?      �?              �?���                      H@      k@      H@      k@      H@      k@                             �p@                        0   G   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           h@        ��                     t� t                         �?      �?              �?���                      R@      k@      R@      k@      R@      k@                             �p@                        H   _   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           h@        ��                     u� t                         �?      �?              �?���                      X@      k@      X@      k@      X@      k@                             �p@                        `   w   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @h@        ��                     v� t                         �?      �?              �?���                      ^@      k@      ^@      k@      ^@      k@                             �p@                        x   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `h@        ��                     w� t                         �?      �?              �?���                      b@      k@      b@      k@      b@      k@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �h@        ��                     x� t                         �?      �?              �?���                      e@      k@      e@      k@      e@      k@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �h@        ��                     y� t                         �?      �?              �?���                      h@      k@      h@      k@      h@      k@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �h@        ��                     z� t                         �?      �?              �?���                      k@      k@      k@      k@      k@      k@                             �p@                        �   �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �h@        ��                     {� t                         �?      �?              �?���                      n@      k@      n@      k@      n@      k@                             �p@                        �     �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           i@        ��                     |� t                         �?      �?              �?���                     �p@      k@     �p@      k@     �p@      k@                             �p@                            �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           i@        ��                     }� t                         �?      �?              �?���                      r@      k@      r@      k@      r@      k@                             �p@                           7  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @i@        ��                     ~� t                         �?      �?              �?���                     �s@      k@     �s@      k@     �s@      k@                             �p@                        8  O  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `i@        ��                     � t                         �?      �?              �?���                      u@      k@      u@      k@      u@      k@                             �p@                        P  g  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �i@        ��                     �� t                         �?      �?              �?���                     �v@      k@     �v@      k@     �v@      k@                             �p@                        h    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �i@        ��                     �� t                         �?      �?              �?���                      x@      k@      x@      k@      x@      k@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �i@        ��                     �� t                         �?      �?              �?���                     �y@      k@     �y@      k@     �y@      k@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �i@        ��                     �� t                         �?      �?              �?���                      {@      k@      {@      k@      {@      k@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           j@        ��                     �� t                         �?      �?              �?���                     �|@      k@     �|@      k@     �|@      k@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           j@        ��                     �� t                         �?      �?              �?���                      ~@      k@      ~@      k@      ~@      k@                             �p@                        �  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @j@        ��                     �� t                         �?      �?              �?���                     �@      k@     �@      k@     �@      k@                             �p@                        �    �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `j@        ��                     �� t                         �?      �?              �?���                     ��@      k@     ��@      k@     ��@      k@                             �p@                          '  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �j@        ��                     �� t                         �?      �?              �?���                     @�@      k@     @�@      k@     @�@      k@                             �p@                        (  ?  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �j@        ��                     �� t                         �?      �?              �?���                      �@      k@      �@      k@      �@      k@                             �p@                        @  W  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �j@        ��                     �� t                         �?      �?              �?���                     ��@      k@     ��@      k@     ��@      k@                             �p@                        X  o  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �j@        ��                     �� t          @              �?      �?              �?���                     ��@      k@     ��@      k@     ��@      k@                             �p@                        p  �  �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           k@        ��                     �� t          @              �?      �?              �?���                              n@              n@              n@                             �p@                               �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           k@        ��                     �� t                         �?      �?              �?���                      8@      n@      8@      n@      8@      n@                             �p@                           /   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @k@        ��                     �� t                         �?      �?              �?���                      H@      n@      H@      n@      H@      n@                             �p@                        0   G   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `k@        ��                     �� t                         �?      �?              �?���                      R@      n@      R@      n@      R@      n@                             �p@                        H   _   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �k@        ��                     �� t                         �?      �?              �?���                      X@      n@      X@      n@      X@      n@                             �p@                        `   w   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �k@        ��                     �� t                         �?      �?              �?���                      ^@      n@      ^@      n@      ^@      n@                             �p@                        x   �   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �k@        ��                     �� t                         �?      �?              �?���                      b@      n@      b@      n@      b@      n@                             �p@                        �   �   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �k@        ��                     �� t                         �?      �?              �?���                      e@      n@      e@      n@      e@      n@                             �p@                        �   �   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           l@        ��                     �� t                         �?      �?              �?���                      h@      n@      h@      n@      h@      n@                             �p@                        �   �   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           l@        ��                     �� t                         �?      �?              �?���                      k@      n@      k@      n@      k@      n@                             �p@                        �   �   �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @l@        ��                     �� t                         �?      �?              �?���                      n@      n@      n@      n@      n@      n@                             �p@                        �     �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `l@        ��                     �� t                         �?      �?              �?���                     �p@      n@     �p@      n@     �p@      n@                             �p@                            �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �l@        ��                     �� t                         �?      �?              �?���                      r@      n@      r@      n@      r@      n@                             �p@                           7  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �l@        ��                     �� t                         �?      �?              �?���                     �s@      n@     �s@      n@     �s@      n@                             �p@                        8  O  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �l@        ��                     �� t                         �?      �?              �?���                      u@      n@      u@      n@      u@      n@                             �p@                        P  g  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �l@        ��                     �� t                         �?      �?              �?���                     �v@      n@     �v@      n@     �v@      n@                             �p@                        h    �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           m@        ��                     �� t                         �?      �?              �?���                      x@      n@      x@      n@      x@      n@                             �p@                        �  �  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           m@        ��                     �� t                         �?      �?              �?���                     �y@      n@     �y@      n@     �y@      n@                             �p@                        �  �  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @m@        ��                     �� t                         �?      �?              �?���                      {@      n@      {@      n@      {@      n@                             �p@                        �  �  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `m@        ��                     �� t                         �?      �?              �?���                     �|@      n@     �|@      n@     �|@      n@                             �p@                        �  �  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �m@        ��                     �� t                         �?      �?              �?���                      ~@      n@      ~@      n@      ~@      n@                             �p@                        �  �  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �m@        ��                     �� t                         �?      �?              �?���                     �@      n@     �@      n@     �@      n@                             �p@                        �    �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �m@        ��                     �� t                         �?      �?              �?���                     ��@      n@     ��@      n@     ��@      n@                             �p@                          '  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �m@        ��                     �� t                         �?      �?              �?���                     @�@      n@     @�@      n@     @�@      n@                             �p@                        (  ?  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           n@        ��                     �� t                         �?      �?              �?���                      �@      n@      �@      n@      �@      n@                             �p@                        @  W  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           n@        ��                     �� t                         �?      �?              �?���                     ��@      n@     ��@      n@     ��@      n@                             �p@                        X  o  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @n@        ��                     �� t          @              �?      �?              �?���                     ��@      n@     ��@      n@     ��@      n@                             �p@                        p  �  �                �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `n@        ��                     �� t          @              �?      �?              �?���                             �p@             �p@             �p@                             �p@                                              �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �n@        ��                     �� t                         �?      �?              �?���                      8@     �p@      8@     �p@      8@     �p@                             �p@                           /                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �n@        ��                     �� t                         �?      �?              �?���                      H@     �p@      H@     �p@      H@     �p@                             �p@                        0   G                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �n@        ��                     �� t                         �?      �?              �?���                      R@     �p@      R@     �p@      R@     �p@                             �p@                        H   _                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �n@        ��                     �� t                         �?      �?              �?���                      X@     �p@      X@     �p@      X@     �p@                             �p@                        `   w                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           o@        ��                     �� t                         �?      �?              �?���                      ^@     �p@      ^@     �p@      ^@     �p@                             �p@                        x   �                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           o@        ��                     �� t                         �?      �?              �?���                      b@     �p@      b@     �p@      b@     �p@                             �p@                        �   �                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @o@        ��                     �� t                         �?      �?              �?���                      e@     �p@      e@     �p@      e@     �p@                             �p@                        �   �                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `o@        ��                     �� t                         �?      �?              �?���                      h@     �p@      h@     �p@      h@     �p@                             �p@                        �   �                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �o@        ��                     �� t                         �?      �?              �?���                      k@     �p@      k@     �p@      k@     �p@                             �p@                        �   �                  �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �o@        ��                     �� t                         �?      �?              �?���                      n@     �p@      n@     �p@      n@     �p@                             �p@                        �                    �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �o@        ��                     �� t                         �?      �?              �?���                     �p@     �p@     �p@     �p@     �p@     �p@                             �p@                                           �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �o@        ��                     �� t                         �?      �?              �?���                      r@     �p@      r@     �p@      r@     �p@                             �p@                           7                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           p@        ��                     �� t                         �?      �?              �?���                     �s@     �p@     �s@     �p@     �s@     �p@                             �p@                        8  O                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          p@        ��                     �� t                         �?      �?              �?���                      u@     �p@      u@     �p@      u@     �p@                             �p@                        P  g                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           p@        ��                     �� t                         �?      �?              �?���                     �v@     �p@     �v@     �p@     �v@     �p@                             �p@                        h                   �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0p@        ��                     �� t                         �?      �?              �?���                      x@     �p@      x@     �p@      x@     �p@                             �p@                        �  �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @p@        ��                     �� t                         �?      �?              �?���                     �y@     �p@     �y@     �p@     �y@     �p@                             �p@                        �  �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pp@        ��                     �� t                         �?      �?              �?���                      {@     �p@      {@     �p@      {@     �p@                             �p@                        �  �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `p@        ��                     �� t                         �?      �?              �?���                     �|@     �p@     �|@     �p@     �|@     �p@                             �p@                        �  �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pp@        ��                     �� t                         �?      �?              �?���                      ~@     �p@      ~@     �p@      ~@     �p@                             �p@                        �  �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t                         �?      �?              �?���                     �@     �p@     �@     �p@     �@     �p@                             �p@                        �                   �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t                         �?      �?              �?���                     ��@     �p@     ��@     �p@     ��@     �p@                             �p@                          '                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t                         �?      �?              �?���                     @�@     �p@     @�@     �p@     @�@     �p@                             �p@                        (  ?                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t                         �?      �?              �?���                      �@     �p@      �@     �p@      �@     �p@                             �p@                        @  W                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t                         �?      �?              �?���                     ��@     �p@     ��@     �p@     ��@     �p@                             �p@                        X  o                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t          @              �?      �?              �?���                     ��@     �p@     ��@     �p@     ��@     �p@                             �p@                        p  �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t          @              �?      �?              �?���                              r@              r@              r@                             �p@                                  7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �p@        ��                     �� t                         �?      �?              �?���                      8@      r@      8@      r@      8@      r@                             �p@                           /      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           q@        ��                     �� t                         �?      �?              �?���                      H@      r@      H@      r@      H@      r@                             �p@                        0   G      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          q@        ��                     �� t                         �?      �?              �?���                      R@      r@      R@      r@      R@      r@                             �p@                        H   _      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           q@        ��                     �� t                         �?      �?              �?���                      X@      r@      X@      r@      X@      r@                             �p@                        `   w      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0q@        ��                     �� t                         �?      �?              �?���                      ^@      r@      ^@      r@      ^@      r@                             �p@                        x   �      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @q@        ��                     �� t                         �?      �?              �?���                      b@      r@      b@      r@      b@      r@                             �p@                        �   �      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pq@        ��                     �� t                         �?      �?              �?���                      e@      r@      e@      r@      e@      r@                             �p@                        �   �      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `q@        ��                     �� t                         �?      �?              �?���                      h@      r@      h@      r@      h@      r@                             �p@                        �   �      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pq@        ��                     �� t                         �?      �?              �?���                      k@      r@      k@      r@      k@      r@                             �p@                        �   �      7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                      n@      r@      n@      r@      n@      r@                             �p@                        �        7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                     �p@      r@     �p@      r@     �p@      r@                             �p@                               7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                      r@      r@      r@      r@      r@      r@                             �p@                           7     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                     �s@      r@     �s@      r@     �s@      r@                             �p@                        8  O     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                      u@      r@      u@      r@      u@      r@                             �p@                        P  g     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                     �v@      r@     �v@      r@     �v@      r@                             �p@                        h       7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                      x@      r@      x@      r@      x@      r@                             �p@                        �  �     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �q@        ��                     �� t                         �?      �?              �?���                     �y@      r@     �y@      r@     �y@      r@                             �p@                        �  �     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           r@        ��                     �� t                         �?      �?              �?���                      {@      r@      {@      r@      {@      r@                             �p@                        �  �     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          r@        ��                     �� t                         �?      �?              �?���                     �|@      r@     �|@      r@     �|@      r@                             �p@                        �  �     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           r@        ��                     �� t                         �?      �?              �?���                      ~@      r@      ~@      r@      ~@      r@                             �p@                        �  �     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0r@        ��                     �� t                         �?      �?              �?���                     �@      r@     �@      r@     �@      r@                             �p@                        �       7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @r@        ��                     �� t                         �?      �?              �?���                     ��@      r@     ��@      r@     ��@      r@                             �p@                          '     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pr@        ��                     �� t                         �?      �?              �?���                     @�@      r@     @�@      r@     @�@      r@                             �p@                        (  ?     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `r@        ��                     �� t                         �?      �?              �?���                      �@      r@      �@      r@      �@      r@                             �p@                        @  W     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pr@        ��                     �� t                         �?      �?              �?���                     ��@      r@     ��@      r@     ��@      r@                             �p@                        X  o     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t          @              �?      �?              �?���                     ��@      r@     ��@      r@     ��@      r@                             �p@                        p  �     7             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t          @              �?      �?              �?���                             �s@             �s@             �s@                             �p@                               8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t                         �?      �?              �?���                      8@     �s@      8@     �s@      8@     �s@                             �p@                           /   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t                         �?      �?              �?���                      H@     �s@      H@     �s@      H@     �s@                             �p@                        0   G   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t                         �?      �?              �?���                      R@     �s@      R@     �s@      R@     �s@                             �p@                        H   _   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t                         �?      �?              �?���                      X@     �s@      X@     �s@      X@     �s@                             �p@                        `   w   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t                         �?      �?              �?���                      ^@     �s@      ^@     �s@      ^@     �s@                             �p@                        x   �   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �r@        ��                     �� t                         �?      �?              �?���                      b@     �s@      b@     �s@      b@     �s@                             �p@                        �   �   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           s@        ��                     �� t                         �?      �?              �?���                      e@     �s@      e@     �s@      e@     �s@                             �p@                        �   �   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          s@        ��                     �� t                         �?      �?              �?���                      h@     �s@      h@     �s@      h@     �s@                             �p@                        �   �   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           s@        ��                     �� t                         �?      �?              �?���                      k@     �s@      k@     �s@      k@     �s@                             �p@                        �   �   8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0s@        ��                     �� t                         �?      �?              �?���                      n@     �s@      n@     �s@      n@     �s@                             �p@                        �     8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @s@        ��                     �� t                         �?      �?              �?���                     �p@     �s@     �p@     �s@     �p@     �s@                             �p@                            8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Ps@        ��                     �� t                         �?      �?              �?���                      r@     �s@      r@     �s@      r@     �s@                             �p@                           7  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `s@        ��                     �� t                         �?      �?              �?���                     �s@     �s@     �s@     �s@     �s@     �s@                             �p@                        8  O  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          ps@        ��                     �� t                         �?      �?              �?���                      u@     �s@      u@     �s@      u@     �s@                             �p@                        P  g  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                     �v@     �s@     �v@     �s@     �v@     �s@                             �p@                        h    8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                      x@     �s@      x@     �s@      x@     �s@                             �p@                        �  �  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                     �y@     �s@     �y@     �s@     �y@     �s@                             �p@                        �  �  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                      {@     �s@      {@     �s@      {@     �s@                             �p@                        �  �  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                     �|@     �s@     �|@     �s@     �|@     �s@                             �p@                        �  �  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                      ~@     �s@      ~@     �s@      ~@     �s@                             �p@                        �  �  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                     �@     �s@     �@     �s@     �@     �s@                             �p@                        �    8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �s@        ��                     �� t                         �?      �?              �?���                     ��@     �s@     ��@     �s@     ��@     �s@                             �p@                          '  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           t@        ��                     �� t                         �?      �?              �?���                     @�@     �s@     @�@     �s@     @�@     �s@                             �p@                        (  ?  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          t@        ��                     �� t                         �?      �?              �?���                      �@     �s@      �@     �s@      �@     �s@                             �p@                        @  W  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           t@        ��                     �� t                         �?      �?              �?���                     ��@     �s@     ��@     �s@     ��@     �s@                             �p@                        X  o  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0t@        ��                     �� t          @              �?      �?              �?���                     ��@     �s@     ��@     �s@     ��@     �s@                             �p@                        p  �  8  O             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @t@        ��                     �� t          @              �?      �?              �?���                              u@              u@              u@                             �p@                               P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pt@        ��                     �� t                         �?      �?              �?���                      8@      u@      8@      u@      8@      u@                             �p@                           /   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `t@        ��                     �� t                         �?      �?              �?���                      H@      u@      H@      u@      H@      u@                             �p@                        0   G   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pt@        ��                     �� t                         �?      �?              �?���                      R@      u@      R@      u@      R@      u@                             �p@                        H   _   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                     �� t                         �?      �?              �?���                      X@      u@      X@      u@      X@      u@                             �p@                        `   w   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                     �� t                         �?      �?              �?���                      ^@      u@      ^@      u@      ^@      u@                             �p@                        x   �   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                     �� t                         �?      �?              �?���                      b@      u@      b@      u@      b@      u@                             �p@                        �   �   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                     �� t                         �?      �?              �?���                      e@      u@      e@      u@      e@      u@                             �p@                        �   �   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                      � t                         �?      �?              �?���                      h@      u@      h@      u@      h@      u@                             �p@                        �   �   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                     � t                         �?      �?              �?���                      k@      u@      k@      u@      k@      u@                             �p@                        �   �   P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                     � t                         �?      �?              �?���                      n@      u@      n@      u@      n@      u@                             �p@                        �     P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �t@        ��                     � t                         �?      �?              �?���                     �p@      u@     �p@      u@     �p@      u@                             �p@                            P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           u@        ��                     � t                         �?      �?              �?���                      r@      u@      r@      u@      r@      u@                             �p@                           7  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          u@        ��                     � t                         �?      �?              �?���                     �s@      u@     �s@      u@     �s@      u@                             �p@                        8  O  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           u@        ��                     � t                         �?      �?              �?���                      u@      u@      u@      u@      u@      u@                             �p@                        P  g  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0u@        ��                     � t                         �?      �?              �?���                     �v@      u@     �v@      u@     �v@      u@                             �p@                        h    P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @u@        ��                     � t                         �?      �?              �?���                      x@      u@      x@      u@      x@      u@                             �p@                        �  �  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pu@        ��                     	� t                         �?      �?              �?���                     �y@      u@     �y@      u@     �y@      u@                             �p@                        �  �  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `u@        ��                     
� t                         �?      �?              �?���                      {@      u@      {@      u@      {@      u@                             �p@                        �  �  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pu@        ��                     � t                         �?      �?              �?���                     �|@      u@     �|@      u@     �|@      u@                             �p@                        �  �  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t                         �?      �?              �?���                      ~@      u@      ~@      u@      ~@      u@                             �p@                        �  �  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t                         �?      �?              �?���                     �@      u@     �@      u@     �@      u@                             �p@                        �    P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t                         �?      �?              �?���                     ��@      u@     ��@      u@     ��@      u@                             �p@                          '  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t                         �?      �?              �?���                     @�@      u@     @�@      u@     @�@      u@                             �p@                        (  ?  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t                         �?      �?              �?���                      �@      u@      �@      u@      �@      u@                             �p@                        @  W  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t                         �?      �?              �?���                     ��@      u@     ��@      u@     ��@      u@                             �p@                        X  o  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t          @              �?      �?              �?���                     ��@      u@     ��@      u@     ��@      u@                             �p@                        p  �  P  g             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �u@        ��                     � t          @              �?      �?              �?���                             �v@             �v@             �v@                             �p@                               h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           v@        ��                     � t                         �?      �?              �?���                      8@     �v@      8@     �v@      8@     �v@                             �p@                           /   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          v@        ��                     � t                         �?      �?              �?���                      H@     �v@      H@     �v@      H@     �v@                             �p@                        0   G   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           v@        ��                     � t                         �?      �?              �?���                      R@     �v@      R@     �v@      R@     �v@                             �p@                        H   _   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0v@        ��                     � t                         �?      �?              �?���                      X@     �v@      X@     �v@      X@     �v@                             �p@                        `   w   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @v@        ��                     � t                         �?      �?              �?���                      ^@     �v@      ^@     �v@      ^@     �v@                             �p@                        x   �   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pv@        ��                     � t                         �?      �?              �?���                      b@     �v@      b@     �v@      b@     �v@                             �p@                        �   �   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `v@        ��                     � t                         �?      �?              �?���                      e@     �v@      e@     �v@      e@     �v@                             �p@                        �   �   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pv@        ��                     � t                         �?      �?              �?���                      h@     �v@      h@     �v@      h@     �v@                             �p@                        �   �   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                     � t                         �?      �?              �?���                      k@     �v@      k@     �v@      k@     �v@                             �p@                        �   �   h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                     � t                         �?      �?              �?���                      n@     �v@      n@     �v@      n@     �v@                             �p@                        �     h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                     � t                         �?      �?              �?���                     �p@     �v@     �p@     �v@     �p@     �v@                             �p@                            h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                     � t                         �?      �?              �?���                      r@     �v@      r@     �v@      r@     �v@                             �p@                           7  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                      � t                         �?      �?              �?���                     �s@     �v@     �s@     �v@     �s@     �v@                             �p@                        8  O  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                     !� t                         �?      �?              �?���                      u@     �v@      u@     �v@      u@     �v@                             �p@                        P  g  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                     "� t                         �?      �?              �?���                     �v@     �v@     �v@     �v@     �v@     �v@                             �p@                        h    h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �v@        ��                     #� t                         �?      �?              �?���                      x@     �v@      x@     �v@      x@     �v@                             �p@                        �  �  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           w@        ��                     $� t                         �?      �?              �?���                     �y@     �v@     �y@     �v@     �y@     �v@                             �p@                        �  �  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          w@        ��                     %� t                         �?      �?              �?���                      {@     �v@      {@     �v@      {@     �v@                             �p@                        �  �  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           w@        ��                     &� t                         �?      �?              �?���                     �|@     �v@     �|@     �v@     �|@     �v@                             �p@                        �  �  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0w@        ��                     '� t                         �?      �?              �?���                      ~@     �v@      ~@     �v@      ~@     �v@                             �p@                        �  �  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @w@        ��                     (� t                         �?      �?              �?���                     �@     �v@     �@     �v@     �@     �v@                             �p@                        �    h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pw@        ��                     )� t                         �?      �?              �?���                     ��@     �v@     ��@     �v@     ��@     �v@                             �p@                          '  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `w@        ��                     *� t                         �?      �?              �?���                     @�@     �v@     @�@     �v@     @�@     �v@                             �p@                        (  ?  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pw@        ��                     +� t                         �?      �?              �?���                      �@     �v@      �@     �v@      �@     �v@                             �p@                        @  W  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     ,� t                         �?      �?              �?���                     ��@     �v@     ��@     �v@     ��@     �v@                             �p@                        X  o  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     -� t          @              �?      �?              �?���                     ��@     �v@     ��@     �v@     ��@     �v@                             �p@                        p  �  h               �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     .� t          @              �?      �?              �?���                              x@              x@              x@                             �p@                               �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     /� t                         �?      �?              �?���                      8@      x@      8@      x@      8@      x@                             �p@                           /   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     0� t                         �?      �?              �?���                      H@      x@      H@      x@      H@      x@                             �p@                        0   G   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     1� t                         �?      �?              �?���                      R@      x@      R@      x@      R@      x@                             �p@                        H   _   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     2� t                         �?      �?              �?���                      X@      x@      X@      x@      X@      x@                             �p@                        `   w   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �w@        ��                     3� t                         �?      �?              �?���                      ^@      x@      ^@      x@      ^@      x@                             �p@                        x   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           x@        ��                     4� t                         �?      �?              �?���                      b@      x@      b@      x@      b@      x@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          x@        ��                     5� t                         �?      �?              �?���                      e@      x@      e@      x@      e@      x@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           x@        ��                     6� t                         �?      �?              �?���                      h@      x@      h@      x@      h@      x@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0x@        ��                     7� t                         �?      �?              �?���                      k@      x@      k@      x@      k@      x@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @x@        ��                     8� t                         �?      �?              �?���                      n@      x@      n@      x@      n@      x@                             �p@                        �     �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Px@        ��                     9� t                         �?      �?              �?���                     �p@      x@     �p@      x@     �p@      x@                             �p@                            �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `x@        ��                     :� t                         �?      �?              �?���                      r@      x@      r@      x@      r@      x@                             �p@                           7  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          px@        ��                     ;� t                         �?      �?              �?���                     �s@      x@     �s@      x@     �s@      x@                             �p@                        8  O  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     <� t                         �?      �?              �?���                      u@      x@      u@      x@      u@      x@                             �p@                        P  g  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     =� t                         �?      �?              �?���                     �v@      x@     �v@      x@     �v@      x@                             �p@                        h    �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     >� t                         �?      �?              �?���                      x@      x@      x@      x@      x@      x@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     ?� t                         �?      �?              �?���                     �y@      x@     �y@      x@     �y@      x@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     @� t                         �?      �?              �?���                      {@      x@      {@      x@      {@      x@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     A� t                         �?      �?              �?���                     �|@      x@     �|@      x@     �|@      x@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     B� t                         �?      �?              �?���                      ~@      x@      ~@      x@      ~@      x@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �x@        ��                     C� t                         �?      �?              �?���                     �@      x@     �@      x@     �@      x@                             �p@                        �    �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           y@        ��                     D� t                         �?      �?              �?���                     ��@      x@     ��@      x@     ��@      x@                             �p@                          '  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          y@        ��                     E� t                         �?      �?              �?���                     @�@      x@     @�@      x@     @�@      x@                             �p@                        (  ?  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           y@        ��                     F� t                         �?      �?              �?���                      �@      x@      �@      x@      �@      x@                             �p@                        @  W  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0y@        ��                     G� t                         �?      �?              �?���                     ��@      x@     ��@      x@     ��@      x@                             �p@                        X  o  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @y@        ��                     H� t          @              �?      �?              �?���                     ��@      x@     ��@      x@     ��@      x@                             �p@                        p  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Py@        ��                     I� t          @              �?      �?              �?���                             �y@             �y@             �y@                             �p@                               �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `y@        ��                     J� t          @              �?      �?              �?���                      8@     �y@      8@     �y@      8@     �y@                             �p@                           /   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          py@        ��                     K� t          @              �?      �?              �?���                      H@     �y@      H@     �y@      H@     �y@                             �p@                        0   G   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     L� t          @              �?      �?              �?���                      R@     �y@      R@     �y@      R@     �y@                             �p@                        H   _   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     M� t          @              �?      �?              �?���                      X@     �y@      X@     �y@      X@     �y@                             �p@                        `   w   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     N� t          @              �?      �?              �?���                      ^@     �y@      ^@     �y@      ^@     �y@                             �p@                        x   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     O� t          @              �?      �?              �?���                      b@     �y@      b@     �y@      b@     �y@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     P� t          @              �?      �?              �?���                      e@     �y@      e@     �y@      e@     �y@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     Q� t          @              �?      �?              �?���                      h@     �y@      h@     �y@      h@     �y@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     R� t          @              �?      �?              �?���                      k@     �y@      k@     �y@      k@     �y@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �y@        ��                     S� t          @              �?      �?              �?���                      n@     �y@      n@     �y@      n@     �y@                             �p@                        �     �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           z@        ��                     T� t          @              �?      �?              �?���                     �p@     �y@     �p@     �y@     �p@     �y@                             �p@                            �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          z@        ��                     U� t          @              �?      �?              �?���                      r@     �y@      r@     �y@      r@     �y@                             �p@                           7  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           z@        ��                     V� t          @              �?      �?              �?���                     �s@     �y@     �s@     �y@     �s@     �y@                             �p@                        8  O  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          0z@        ��                     W� t          @              �?      �?              �?���                      u@     �y@      u@     �y@      u@     �y@                             �p@                        P  g  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          @z@        ��                     X� t          @              �?      �?              �?���                     �v@     �y@     �v@     �y@     �v@     �y@                             �p@                        h    �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          Pz@        ��                     Y� t          @              �?      �?              �?���                      x@     �y@      x@     �y@      x@     �y@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          `z@        ��                     Z� t          @              �?      �?              �?���                     �y@     �y@     �y@     �y@     �y@     �y@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          pz@        ��                     [� t          @              �?      �?              �?���                      {@     �y@      {@     �y@      {@     �y@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     \� t          @              �?      �?              �?���                     �|@     �y@     �|@     �y@     �|@     �y@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     ]� t          @              �?      �?              �?���                      ~@     �y@      ~@     �y@      ~@     �y@                             �p@                        �  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     ^� t          @              �?      �?              �?���                     �@     �y@     �@     �y@     �@     �y@                             �p@                        �    �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     _� t          @              �?      �?              �?���                     ��@     �y@     ��@     �y@     ��@     �y@                             �p@                          '  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     `� t          @              �?      �?              �?���                     @�@     �y@     @�@     �y@     @�@     �y@                             �p@                        (  ?  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     a� t          @              �?      �?              �?���                      �@     �y@      �@     �y@      �@     �y@                             �p@                        @  W  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     b� t          @              �?      �?              �?���                     ��@     �y@     ��@     �y@     ��@     �y@                             �p@                        X  o  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��          �z@        ��                     c� t          @              �?      �?              �?���                     ��@     �y@     ��@     �y@     ��@     �y@                             �p@                        p  �  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ��           {@        ��                     �� �                 �?      �?      �?              �?��� ����                 X@      {@      X@      {@      X@      {@                             �p@                        `   w   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����                 n@      {@      n@      {@      n@      {@                             �p@                        �     �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����                 k@      {@      k@      {@      k@      {@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����                 r@      {@      r@      {@      r@      {@                             �p@                           7  �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����                 H@      {@      H@      {@      H@      {@                             �p@                        (   O   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����                 ^@      {@      ^@      {@      ^@      {@                             �p@                        x   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �     ш            	   basic.lef    �� �                 �?      �?      �?              �?��� ����                 b@      {@      b@      {@      b@      {@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����                 e@      {@      e@      {@      e@      {@                             �p@                        �   �   �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� 
                 �?      �?      �?              �?���                     ��@      8@     ��@      8@     ��@      8@                             �p@                        X  o     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                  �?      �?      �?              �?���                      �@      8@      �@      8@      �@      8@                             �p@                        @  W     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                          �?      �?              �?���                     @�@      8@     @�@      8@     @�@      8@                             �p@                        (  ?     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� '                 �?      �?      �?              �?���                     �@      8@     �@      8@     �@      8@                             �p@                        �       /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                          �?      �?              �?���                      {@      8@      {@      8@      {@      8@                             �p@                        �  �     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                  �?      �?      �?              �?���                     �y@      8@     �y@      8@     �y@      8@                             �p@                        �  �     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?���                      ~@      8@      ~@      8@      ~@      8@                             �p@                        �  �     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� E                 �?      �?      �?              �?���                     �|@      8@     �|@      8@     �|@      8@                             �p@                        �  �     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� N                 �?      �?      �?              �?���                      x@      8@      x@      8@      x@      8@                             �p@                        �  �     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                  �?      �?      �?              �?���                     �v@      8@     �v@      8@     �v@      8@                             �p@                        h       /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                  �?      �?      �?              �?���                      u@      8@      u@      8@      u@      8@                             �p@                        P  g     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                  �?      �?      �?              �?���                     ��@      8@     ��@      8@     ��@      8@                             �p@                          '     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����                �p@      {@     �p@      {@     �p@      {@                             �p@                            �  �             �   ������������������������������������������������        ����                              �?                            ����              �?    �      ��                          �?      �?              �?���                     ��@      8@     ��@      8@     ��@      8@                             �p@                        p  �     /              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� ����     X�@      �?      �?      �?              �?��� ����                  H@              H@              H@                                     �p@                        `y��`y��`y��`y��             ������������������������������������������������        ����                              �?                            ����              �?    �      �� �                 �?      �?      �?              �?��� ����      �                 h@              h@              h@                             �p@                           �   �   �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      d� t         �?              �?      �?              �?���            �         8@      k@     �|@      n@      8@      k@                             �p@                           /   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      e� t          @              �?      �?              �?���            �         H@      k@      ~@      n@      H@      k@                             �p@                        0   G   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      f� t         @              �?      �?              �?���            �         R@      k@     �@      n@      R@      k@                             �p@                        H   _   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      g� t         @              �?      �?              �?���            �         X@      k@     ��@      n@      X@      k@                             �p@                        `   w   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      h� t         @              �?      �?              �?���            �         ^@      k@     @�@      n@      ^@      k@                             �p@                        x   �   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      i� t         @              �?      �?              �?���            �         b@      k@      �@      n@      b@      k@                             �p@                        �   �   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      j� t         @              �?      �?              �?���            �         e@      k@     ��@      n@      e@      k@                             �p@                        �   �   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      k� t          @              �?      �?              �?���            �         h@      k@     ��@      n@      h@      k@                             �p@                        �   �   �   �               �   ������������������������������������������������        ����                              �?                            ����              �?    �      l� t         "@              �?      �?              �?���            �         8@      n@     �|@     �p@      8@      n@                             �p@                           /   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      m� t         $@              �?      �?              �?���            �         H@      n@      ~@     �p@      H@      n@                             �p@                        0   G   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      n� t         &@              �?      �?              �?���            �         R@      n@     �@     �p@      R@      n@                             �p@                        H   _   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      o� t         (@              �?      �?              �?���            �         X@      n@     ��@     �p@      X@      n@                             �p@                        `   w   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      p� t         *@              �?      �?              �?���            �         ^@      n@     @�@     �p@      ^@      n@                             �p@                        x   �   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      q� t         ,@              �?      �?              �?���            �         b@      n@      �@     �p@      b@      n@                             �p@                        �   �   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      r� t         .@              �?      �?              �?���            �         e@      n@     ��@     �p@      e@      n@                             �p@                        �   �   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      s� t         0@              �?      �?              �?���            �         h@      n@     ��@     �p@      h@      n@                             �p@                        �   �   �                 �   ������������������������������������������������        ����                              �?                            ����              �?    �      t� t         1@              �?      �?              �?���            �         8@     �p@     �|@      r@      8@     �p@                             �p@                           /                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      u� t         2@              �?      �?              �?���            �         H@     �p@      ~@      r@      H@     �p@                             �p@                        0   G                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      v� t         3@              �?      �?              �?���            �         R@     �p@     �@      r@      R@     �p@                             �p@                        H   _                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      w� t         4@              �?      �?              �?���            �         X@     �p@     ��@      r@      X@     �p@                             �p@                        `   w                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      x� t         5@              �?      �?              �?���            �         ^@     �p@     @�@      r@      ^@     �p@                             �p@                        x   �                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      y� t         6@              �?      �?              �?���            �         b@     �p@      �@      r@      b@     �p@                             �p@                        �   �                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      z� t         7@              �?      �?              �?���            �         e@     �p@     ��@      r@      e@     �p@                             �p@                        �   �                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      {� t         8@              �?      �?              �?���            �         h@     �p@     ��@      r@      h@     �p@                             �p@                        �   �                   �   ������������������������������������������������        ����                              �?                            ����              �?    �      |� t         9@              �?      �?              �?���            �         8@      r@     �|@     �s@      8@      r@                             �p@                           /      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      }� t         :@              �?      �?              �?���            �         H@      r@      ~@     �s@      H@      r@                             �p@                        0   G      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      ~� t         ;@              �?      �?              �?���            �         R@      r@     �@     �s@      R@      r@                             �p@                        H   _      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      � t         <@              �?      �?              �?���            �         X@      r@     ��@     �s@      X@      r@                             �p@                        `   w      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         =@              �?      �?              �?���            �         ^@      r@     @�@     �s@      ^@      r@                             �p@                        x   �      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         >@              �?      �?              �?���            �         b@      r@      �@     �s@      b@      r@                             �p@                        �   �      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         ?@              �?      �?              �?���            �         e@      r@     ��@     �s@      e@      r@                             �p@                        �   �      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         @@              �?      �?              �?���            �         h@      r@     ��@     �s@      h@      r@                             �p@                        �   �      7              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �@@              �?      �?              �?���            �         8@     �s@     �|@      u@      8@     �s@                             �p@                           /   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         A@              �?      �?              �?���            �         H@     �s@      ~@      u@      H@     �s@                             �p@                        0   G   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �A@              �?      �?              �?���            �         R@     �s@     �@      u@      R@     �s@                             �p@                        H   _   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         B@              �?      �?              �?���            �         X@     �s@     ��@      u@      X@     �s@                             �p@                        `   w   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �B@              �?      �?              �?���            �         ^@     �s@     @�@      u@      ^@     �s@                             �p@                        x   �   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         C@              �?      �?              �?���            �         b@     �s@      �@      u@      b@     �s@                             �p@                        �   �   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �C@              �?      �?              �?���            �         e@     �s@     ��@      u@      e@     �s@                             �p@                        �   �   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         D@              �?      �?              �?���            �         h@     �s@     ��@      u@      h@     �s@                             �p@                        �   �   8  O              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �D@              �?      �?              �?���            �         8@      u@     �|@     �v@      8@      u@                             �p@                           /   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         E@              �?      �?              �?���            �         H@      u@      ~@     �v@      H@      u@                             �p@                        0   G   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �E@              �?      �?              �?���            �         R@      u@     �@     �v@      R@      u@                             �p@                        H   _   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         F@              �?      �?              �?���            �         X@      u@     ��@     �v@      X@      u@                             �p@                        `   w   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �F@              �?      �?              �?���            �         ^@      u@     @�@     �v@      ^@      u@                             �p@                        x   �   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         G@              �?      �?              �?���            �         b@      u@      �@     �v@      b@      u@                             �p@                        �   �   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �G@              �?      �?              �?���            �         e@      u@     ��@     �v@      e@      u@                             �p@                        �   �   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         H@              �?      �?              �?���            �         h@      u@     ��@     �v@      h@      u@                             �p@                        �   �   P  g              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �H@              �?      �?              �?���            �         8@     �v@     �|@      x@      8@     �v@                             �p@                           /   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         I@              �?      �?              �?���            �         H@     �v@      ~@      x@      H@     �v@                             �p@                        0   G   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �I@              �?      �?              �?���            �         R@     �v@     �@      x@      R@     �v@                             �p@                        H   _   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         J@              �?      �?              �?���            �         X@     �v@     ��@      x@      X@     �v@                             �p@                        `   w   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �J@              �?      �?              �?���            �         ^@     �v@     @�@      x@      ^@     �v@                             �p@                        x   �   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         K@              �?      �?              �?���            �         b@     �v@      �@      x@      b@     �v@                             �p@                        �   �   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �K@              �?      �?              �?���            �         e@     �v@     ��@      x@      e@     �v@                             �p@                        �   �   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         L@              �?      �?              �?���            �         h@     �v@     ��@      x@      h@     �v@                             �p@                        �   �   h                �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �L@              �?      �?              �?���            �         8@      x@     �|@     �y@      8@      x@                             �p@                           /   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         M@              �?      �?              �?���            �         H@      x@      ~@     �y@      H@      x@                             �p@                        0   G   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �M@              �?      �?              �?���            �         R@      x@     �@     �y@      R@      x@                             �p@                        H   _   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         N@              �?      �?              �?���            �         X@      x@     ��@     �y@      X@      x@                             �p@                        `   w   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �N@              �?      �?              �?���            �         ^@      x@     @�@     �y@      ^@      x@                             �p@                        x   �   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         O@              �?      �?              �?���            �         b@      x@      �@     �y@      b@      x@                             �p@                        �   �   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t        �O@              �?      �?              �?���            �         e@      x@     ��@     �y@      e@      x@                             �p@                        �   �   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �� t         P@              �?      �?              �?���            �         h@      x@     ��@     �y@      h@      x@                             �p@                        �   �   �  �              �   ������������������������������������������������        ����                              �?                            ����              �?    �      �O [                 �?      �?      �?              �?��� ����     �V�                                 k@                                             �p@                            �      .              G   ������������������������������������������������        ����                              �?                            ����              �?    �     Ĉ           �?        �O \                 �?      �?      �?              �?��� ����     �V�                 {@              n@              {@                             �p@                            �  �  �             H   ������������������������������������������������        ����                              �?                            ����              �?    �     Ĉ           �?        �� ����     X�@      �?      �?      �?              �?��� ����      Y�          8@              8@              8@                                     �p@                        `y��`y��`y��`y��           F   ������������������������������������������������        ����                              �?                            ����              �?    �     ��               Custom Levels    ��                                        È               Level Editor                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �O �� 